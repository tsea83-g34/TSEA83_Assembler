mem := (
--$PROGRAM
X"move r13 r15: cfdf0000",
X"load r0 r13 2 [2]: 810d0002",
X"cmpi r0 1: e3000001",
X"breq L0: 1b000003",
X"addi r0 r14 0: 8b0e0000",
X"rjmp L1: 33000002",
X"addi r0 r14 1: 8b0e0001",
X"cmpi r0 1: e3000001",
X"brne L2: 1f000006",
X"addi r12 r14 1: 8bce0001",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 13: 8fdd000d",
X"rjmprg r13: efd00000",
X"load r1 r13 2 [2]: 811d0002",
X"cmpi r1 2: e3020002",
X"breq L3: 1b000003",
X"addi r1 r14 0: 8b1e0000",
X"rjmp L4: 33000002",
X"addi r1 r14 1: 8b1e0001",
X"cmpi r1 1: e3020001",
X"brne L5: 1f000006",
X"addi r12 r14 1: 8bce0001",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 26: 8fdd001a",
X"rjmprg r13: efd00000",
X"subi r15 r15 2: 8fff0002",
X"addi r2 r14 1: 8b2e0001",
X"subi r15 r15 2: 8fff0002",
X"addi r3 r14 1: 8b3e0001",
X"subi r15 r15 2: 8fff0002",
X"addi r4 r14 0: 8b4e0000",
X"subi r15 r15 2: 8fff0002",
X"addi r5 r14 2: 8b5e0002",
X"store r13 r2 -2 [2]: d1d2fffe",
X"store r13 r3 -4 [2]: d1d3fffc",
X"store r13 r4 -6 [2]: d1d4fffa",
X"store r13 r5 -8 [2]: d1d5fff8",
X"load r0 r13 -8 [2]: 810dfff8",
X"load r1 r13 2 [2]: 811d0002",
X"cmp r0 r1: df002000",
X"brne L8: 1f000003",
X"addi r0 r14 0: 8b0e0000",
X"rjmp L9: 33000002",
X"addi r0 r14 1: 8b0e0001",
X"cmpi r0 1: e3000001",
X"brne L7: 1f00001f",
X"load r2 r13 -6 [2]: 812dfffa",
X"cmpi r2 0: e3040000",
X"breq L10: 1b000003",
X"addi r2 r14 0: 8b2e0000",
X"rjmp L11: 33000002",
X"addi r2 r14 1: 8b2e0001",
X"cmpi r2 1: e3040001",
X"brne L12: 1f000006",
X"load r3 r13 -2 [2]: 813dfffe",
X"load r4 r13 -4 [2]: 814dfffc",
X"add r3 r3 r4: 93334000",
X"move r5 r3: cf530000",
X"addi r6 r14 1: 8b6e0001",
X"cmpi r6 1: e30c0001",
X"breq L13: 1b000003",
X"addi r6 r14 0: 8b6e0000",
X"rjmp L14: 33000002",
X"addi r6 r14 1: 8b6e0001",
X"cmpi r6 1: e30c0001",
X"brne L15: 1f000004",
X"add r4 r4 r5: 93445000",
X"move r3 r4: cf340000",
X"addi r6 r14 0: 8b6e0000",
X"addi r1 r1 1: 8b110001",
X"move r4 r1: cf410000",
X"store r13 r3 -4 [2]: d1d3fffc",
X"store r13 r4 2 [2]: d1d40002",
X"store r13 r5 -2 [2]: d1d5fffe",
X"store r13 r6 -6 [2]: d1d6fffa",
X"rjmp L6: 3300ffda",
X"load r0 r13 -6 [2]: 810dfffa",
X"cmpi r0 0: e3000000",
X"breq L16: 1b000003",
X"addi r0 r14 0: 8b0e0000",
X"rjmp L17: 33000002",
X"addi r0 r14 1: 8b0e0001",
X"cmpi r0 1: e3000001",
X"brne L18: 1f000008",
X"load r1 r13 -4 [2]: 811dfffc",
X"move r12 r1: cfc10000",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 92: 8fdd005c",
X"rjmprg r13: efd00000",
X"load r2 r13 -6 [2]: 812dfffa",
X"cmpi r2 1: e3040001",
X"breq L19: 1b000003",
X"addi r2 r14 0: 8b2e0000",
X"rjmp L20: 33000002",
X"addi r2 r14 1: 8b2e0001",
X"cmpi r2 1: e3040001",
X"brne L21: 1f000008",
X"load r3 r13 -2 [2]: 813dfffe",
X"move r12 r3: cfc30000",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 107: 8fdd006b",
X"rjmprg r13: efd00000",
X"addi r15 r15 8: 8bff0008",
X"move r12 r14: cfce0000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 113: 8fdd0071",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"subi r15 r15 2: 8fff0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"addi r0 r14 10: 8b0e000a",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r0 0 [2]: d1f00000",
X"movlo r13 126: f7d0007e",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp fibonacci: 3300ff83",
X"addi r15 r15 4: 8bff0004",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"move r0 r12: cf0c0000",
X"addi r12 r14 0: 8bce0000",
X"addi r15 r15 2: 8bff0002",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 135: 8fdd0087",
X"rjmprg r13: efd00000",
--$PROGRAM_END
others => X"00000000"
);