mem := (
--$DATA
X"68",
X"65",
X"6c",
X"6c",
X"6f",
X"00",
X"ff",
X"aa",
X"aa",
X"dc",
X"fe",
X"34",
X"12",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"fd",
--$DATA_END
others => X"00"
)