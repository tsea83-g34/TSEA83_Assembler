mem := (
--$PROGRAM
"10010011000000000001000000000000",
"10001011000100010000000000000001",
"00001011110100000000000000000000",
"11101111110100000000000000000000",
"00111111110101110000000000000111",
"11011011110100000000000000000000",
"00110011000000001111111111111011",
--$PROGRAM_END
others => X"00000000"
);