mem := (
--$PROGRAM
X"cb001000",
X"c7110001",
X"0b900000",
X"07900000",
X"17980008",
X"db900000",
X"0700fffb",
--$PROGRAM_END
others => X"00000000"
);