mem := (
--$PROGRAM
X"93001000",
X"8b110001",
X"0bd00000",
X"07d00000",
X"17d70007",
X"dbd00000",
X"0700fffb",
--$PROGRAM_END
others => X"00000000"
);