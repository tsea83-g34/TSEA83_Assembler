mem := (
--$DATA

--$DATA_END
others => X"00"
)