mem1 := (
--$DATA1
X"00",
--$DATA1_END
others => X"00"
)

mem2 := (
--$DATA2
X"10",
--$DATA2_END
others => X"00"
)

mem3 := (
--$DATA3

--$DATA3_END
others => X"00"
)

mem4 := (
--$DATA4

--$DATA4_END
others => X"00"
)