mem := (
--$PROGRAM
X"load r0 r14 2 [2]: 810e0002",
X"load r1 r14 4 [2]: 811e0004",
X"mul r0 r0 r1: a7001000",
X"store r14 r0 6 [2]: d1e00006",
X"load r0 r14 6 [2]: 810e0006",
X"store r14 r0 8 [2]: d1e00008",
X"load r0 r14 6 [2]: 810e0006",
X"load r2 r14 10 [2]: 812e000a",
X"add r0 r0 r2: 93002000",
X"store r14 r0 12 [2]: d1e0000c",
X"move r13 r15: cfdf0000",
X"load r0 r13 2 [2]: 810d0002",
X"subi r15 r15 4: 8fff0004",
X"load r1 r13 -4 [4]: 831dfffc",
X"in r1 r0: 0f100000",
X"move r12 r1: cfc10000",
X"addi r15 r15 4: 8bff0004",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 20: 8fdd0014",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"load r0 r13 4 [4]: 830d0004",
X"load r1 r13 10 [2]: 811d000a",
X"out r1 r0: e7100000",
X"move r12 r14: cfce0000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 29: 8fdd001d",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"load r0 r13 4 [4]: 830d0004",
X"load r1 r13 10 [2]: 811d000a",
X"vgaw r1 r0: eb100000",
X"move r12 r14: cfce0000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 38: 8fdd0026",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"load r0 r13 2 [2]: 810d0002",
X"load r1 r13 4 [2]: 811d0004",
X"load r2 r13 6 [2]: 812d0006",
X"cmp r0 r2: df004000",
X"brge L0: 2f000003",
X"addi r0 r14 0: 8b0e0000",
X"rjmp L1: 33000002",
X"addi r0 r14 1: 8b0e0001",
X"load r3 r13 2 [2]: 813d0002",
X"cmp r3 r1: df062000",
X"brlt L2: 23000003",
X"addi r3 r14 0: 8b3e0000",
X"rjmp L3: 33000002",
X"addi r3 r14 1: 8b3e0001",
X"or r0 r0 r3: c3003000",
X"move r12 r0: cfc00000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 59: 8fdd003b",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"load r0 r13 4 [2]: 810d0004",
X"load r1 r13 6 [2]: 811d0006",
X"subi r15 r15 2: 8fff0002",
X"subi r15 r15 2: 8fff0002",
X"addi r2 r14 0: 8b2e0000",
X"store r13 r0 -2 [2]: d1d0fffe",
X"store r13 r2 -4 [2]: d1d2fffc",
X"load r0 r13 -2 [2]: 810dfffe",
X"load r1 r13 6 [2]: 811d0006",
X"cmp r0 r1: df002000",
X"brgt L6: 27000003",
X"addi r0 r14 0: 8b0e0000",
X"rjmp L7: 33000002",
X"addi r0 r14 1: 8b0e0001",
X"cmpi r0 1: e3000001",
X"brne L5: 1f000008",
X"load r2 r13 -2 [2]: 812dfffe",
X"sub r2 r2 r1: 97221000",
X"move r3 r2: cf320000",
X"load r4 r13 -4 [2]: 814dfffc",
X"addi r4 r4 1: 8b440001",
X"move r5 r4: cf540000",
X"rjmp L4: 3300fff1",
X"subi r15 r15 4: 8fff0004",
X"load r0 r13 -4 [2]: 810dfffc",
X"store r13 r0 -8 [4]: d3d0fff8",
X"load r1 r13 -2 [2]: 811dfffe",
X"add r0 r0 r1: 93001000",
X"move r2 r0: cf200000",
X"move r12 r2: cfc20000",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 95: 8fdd005f",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"load r0 r13 4 [4]: 830d0004",
X"load r3 r13 10 [2]: 813d000a",
X"load r4 r14 6 [2]: 814e0006",
X"cmp r3 r4: df068000",
X"brge L8: 2f000003",
X"addi r3 r14 0: 8b3e0000",
X"rjmp L9: 33000002",
X"addi r3 r14 1: 8b3e0001",
X"cmpi r3 1: e3060001",
X"brne L10: 1f000007",
X"addi r12 r14 0: 8bce0000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 111: 8fdd006f",
X"rjmprg r13: efd00000",
X"rjmp L11: 33000001",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r0 r13 10 [2]: 810d000a",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r0 0 [2]: d1f00000",
X"load r1 r13 4 [4]: 831d0004",
X"subi r15 r15 2: 8fff0002",
X"addi r15 r15 -4: 8bfffffc",
X"store r15 r1 0 [4]: d3f10000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 128: f7d00080",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp vga_write: 3300ff9f",
X"addi r15 r15 12: 8bff000c",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r12 r14 1: 8bce0001",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 135: 8fdd0087",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"load r0 r13 4 [4]: 830d0004",
X"load r1 r13 8 [2]: 811d0008",
X"load r2 r13 10 [2]: 812d000a",
X"load r3 r14 14 [2]: 813e000e",
X"cmp r1 r3: df026000",
X"brge L12: 2f000003",
X"addi r1 r14 0: 8b1e0000",
X"rjmp L13: 33000002",
X"addi r1 r14 1: 8b1e0001",
X"load r4 r14 16 [2]: 814e0010",
X"cmp r2 r4: df048000",
X"brge L14: 2f000003",
X"addi r2 r14 0: 8b2e0000",
X"rjmp L15: 33000002",
X"addi r2 r14 1: 8b2e0001",
X"or r1 r1 r2: c3112000",
X"cmpi r1 1: e3020001",
X"brne L16: 1f000007",
X"addi r12 r14 0: 8bce0000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 159: 8fdd009f",
X"rjmprg r13: efd00000",
X"rjmp L17: 33000001",
X"subi r15 r15 2: 8fff0002",
X"load r0 r13 8 [2]: 810d0008",
X"load r1 r14 14 [2]: 811e000e",
X"load r2 r13 10 [2]: 812d000a",
X"mul r1 r1 r2: a7112000",
X"add r0 r0 r1: 93001000",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r0 0 [2]: d1f00000",
X"load r3 r13 4 [4]: 833d0004",
X"subi r15 r15 2: 8fff0002",
X"addi r15 r15 -4: 8bfffffc",
X"store r15 r3 0 [4]: d3f30000",
X"store r13 r0 -2 [2]: d1d0fffe",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 181: f7d000b5",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp vga_write: 3300ff6a",
X"addi r15 r15 10: 8bff000a",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r12 r14 1: 8bce0001",
X"addi r15 r15 2: 8bff0002",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 189: 8fdd00bd",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"load r0 r13 4 [2]: 810d0004",
X"load r1 r13 6 [1]: 801d0006",
X"load r2 r13 7 [1]: 802d0007",
X"load r3 r14 10 [2]: 813e000a",
X"cmp r0 r3: df006000",
X"brge L18: 2f000003",
X"addi r0 r14 0: 8b0e0000",
X"rjmp L19: 33000002",
X"addi r0 r14 1: 8b0e0001",
X"cmpi r0 1: e3000001",
X"brne L20: 1f000007",
X"addi r12 r14 0: 8bce0000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 206: 8fdd00ce",
X"rjmprg r13: efd00000",
X"rjmp L21: 33000001",
X"subi r15 r15 2: 8fff0002",
X"load r0 r14 8 [2]: 810e0008",
X"load r1 r13 4 [2]: 811d0004",
X"add r0 r0 r1: 93001000",
X"subi r15 r15 6: 8fff0006",
X"load r2 r13 6 [1]: 802d0006",
X"store r13 r2 -8 [4]: d3d2fff8",
X"load r3 r13 7 [1]: 803d0007",
X"add r2 r2 r3: 93223000",
X"move r4 r2: cf420000",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r0 0 [2]: d1f00000",
X"subi r15 r15 2: 8fff0002",
X"addi r15 r15 -4: 8bfffffc",
X"store r15 r4 0 [4]: d3f40000",
X"store r13 r0 -2 [2]: d1d0fffe",
X"store r13 r4 -8 [4]: d3d4fff8",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 233: f7d000e9",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp vga_write: 3300ff36",
X"addi r15 r15 12: 8bff000c",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r12 r14 1: 8bce0001",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 241: 8fdd00f1",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"load r0 r13 2 [1]: 800d0002",
X"load r1 r13 3 [1]: 801d0003",
X"load r2 r14 2 [2]: 812e0002",
X"cmp r0 r2: df004000",
X"brge L22: 2f000003",
X"addi r0 r14 0: 8b0e0000",
X"rjmp L23: 33000002",
X"addi r0 r14 1: 8b0e0001",
X"load r3 r14 4 [2]: 813e0004",
X"cmp r1 r3: df026000",
X"brge L24: 2f000003",
X"addi r1 r14 0: 8b1e0000",
X"rjmp L25: 33000002",
X"addi r1 r14 1: 8b1e0001",
X"or r0 r0 r1: c3001000",
X"cmpi r0 1: e3000001",
X"brne L26: 1f000007",
X"addi r12 r14 0: 8bce0000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 264: 8fdd0108",
X"rjmprg r13: efd00000",
X"rjmp L27: 33000001",
X"load r0 r13 2 [1]: 800d0002",
X"move r1 r0: cf100000",
X"load r2 r13 3 [1]: 802d0003",
X"move r3 r2: cf320000",
X"add r0 r0 r2: 93002000",
X"load r4 r14 2 [2]: 814e0002",
X"mul r0 r0 r4: a7004000",
X"move r5 r0: cf500000",
X"addi r12 r14 1: 8bce0001",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 278: 8fdd0116",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"load r0 r14 20 [2]: 810e0014",
X"addi r0 r0 1: 8b000001",
X"move r1 r0: cf100000",
X"store r14 r1 20 [2]: d1e10014",
X"load r2 r14 6 [2]: 812e0006",
X"cmp r1 r2: df024000",
X"brlt L28: 23000003",
X"addi r1 r14 0: 8b1e0000",
X"rjmp L29: 33000002",
X"addi r1 r14 1: 8b1e0001",
X"cmpi r1 1: e3020001",
X"brne L30: 1f000015",
X"load r0 r14 22 [2]: 810e0016",
X"addi r0 r0 1: 8b000001",
X"move r1 r0: cf100000",
X"store r14 r1 22 [2]: d1e10016",
X"load r2 r14 2 [2]: 812e0002",
X"cmp r1 r2: df024000",
X"brge L32: 2f000003",
X"addi r1 r14 0: 8b1e0000",
X"rjmp L33: 33000002",
X"addi r1 r14 1: 8b1e0001",
X"cmpi r1 1: e3020001",
X"brne L34: 1f000008",
X"addi r0 r14 0: 8b0e0000",
X"load r1 r14 24 [2]: 811e0018",
X"addi r1 r1 1: 8b110001",
X"move r2 r1: cf210000",
X"store r14 r0 22 [2]: d1e00016",
X"store r14 r2 24 [2]: d1e20018",
X"rjmp L35: 33000001",
X"rjmp L31: 33000007",
X"addi r0 r14 0: 8b0e0000",
X"addi r1 r14 0: 8b1e0000",
X"addi r2 r14 0: 8b2e0000",
X"store r14 r0 20 [2]: d1e00014",
X"store r14 r1 22 [2]: d1e10016",
X"store r14 r2 24 [2]: d1e20018",
X"move r12 r14: cfce0000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 322: 8fdd0142",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"load r0 r14 20 [2]: 810e0014",
X"subi r0 r0 1: 8f000001",
X"move r1 r0: cf100000",
X"store r14 r1 20 [2]: d1e10014",
X"load r2 r14 6 [2]: 812e0006",
X"cmp r1 r2: df024000",
X"brlt L36: 23000003",
X"addi r1 r14 0: 8b1e0000",
X"rjmp L37: 33000002",
X"addi r1 r14 1: 8b1e0001",
X"cmpi r1 1: e3020001",
X"brne L38: 1f000014",
X"load r0 r14 22 [2]: 810e0016",
X"subi r0 r0 1: 8f000001",
X"move r1 r0: cf100000",
X"store r14 r1 22 [2]: d1e10016",
X"cmpi r1 0: e3020000",
X"brlt L40: 23000003",
X"addi r1 r14 0: 8b1e0000",
X"rjmp L41: 33000002",
X"addi r1 r14 1: 8b1e0001",
X"cmpi r1 1: e3020001",
X"brne L42: 1f000008",
X"addi r0 r14 0: 8b0e0000",
X"load r1 r14 24 [2]: 811e0018",
X"subi r1 r1 1: 8f110001",
X"move r2 r1: cf210000",
X"store r14 r0 22 [2]: d1e00016",
X"store r14 r2 24 [2]: d1e20018",
X"rjmp L43: 33000001",
X"rjmp L39: 3300000b",
X"load r0 r14 6 [2]: 810e0006",
X"subi r0 r0 1: 8f000001",
X"move r1 r0: cf100000",
X"load r2 r14 2 [2]: 812e0002",
X"move r3 r2: cf320000",
X"load r4 r14 4 [2]: 814e0004",
X"move r5 r4: cf540000",
X"store r14 r1 20 [2]: d1e10014",
X"store r14 r3 22 [2]: d1e30016",
X"store r14 r5 24 [2]: d1e50018",
X"move r12 r14: cfce0000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 369: 8fdd0171",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"load r0 r13 2 [2]: 810d0002",
X"load r1 r14 6 [2]: 811e0006",
X"cmp r0 r1: df002000",
X"brge L44: 2f000003",
X"addi r0 r14 0: 8b0e0000",
X"rjmp L45: 33000002",
X"addi r0 r14 1: 8b0e0001",
X"cmpi r0 1: e3000001",
X"brne L46: 1f000007",
X"addi r12 r14 0: 8bce0000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 384: 8fdd0180",
X"rjmprg r13: efd00000",
X"rjmp L47: 33000001",
X"load r0 r14 20 [2]: 810e0014",
X"load r1 r13 2 [2]: 811d0002",
X"add r0 r0 r1: 93001000",
X"move r2 r0: cf200000",
X"store r14 r2 20 [2]: d1e20014",
X"load r3 r14 6 [2]: 813e0006",
X"cmp r2 r3: df046000",
X"brge L48: 2f000003",
X"addi r2 r14 0: 8b2e0000",
X"rjmp L49: 33000002",
X"addi r2 r14 1: 8b2e0001",
X"cmpi r2 1: e3040001",
X"brne L50: 1f000007",
X"load r0 r14 20 [2]: 810e0014",
X"load r1 r14 6 [2]: 811e0006",
X"sub r0 r0 r1: 97001000",
X"move r2 r0: cf200000",
X"store r14 r2 20 [2]: d1e20014",
X"rjmp L51: 33000001",
X"subi r15 r15 4: 8fff0004",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r0 r14 2 [2]: 810e0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r0 0 [2]: d1f00000",
X"load r1 r14 20 [2]: 811e0014",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r1 0 [2]: d1f10000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 420: f7d001a4",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp divide: 3300fe99",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"move r0 r12: cf0c0000",
X"subi r15 r15 4: 8fff0004",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r1 r14 4 [2]: 811e0004",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r1 0 [2]: d1f10000",
X"load r2 r14 20 [2]: 812e0014",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r2 0 [2]: d1f20000",
X"store r13 r0 -4 [4]: d3d0fffc",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 440: f7d001b8",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp divide: 3300fe85",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"move r0 r12: cf0c0000",
X"addi r12 r14 1: 8bce0001",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 449: 8fdd01c1",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"load r0 r14 24 [2]: 810e0018",
X"addi r0 r0 1: 8b000001",
X"move r1 r0: cf100000",
X"store r14 r1 24 [2]: d1e10018",
X"load r2 r14 4 [2]: 812e0004",
X"cmp r1 r2: df024000",
X"brlt L52: 23000003",
X"addi r1 r14 0: 8b1e0000",
X"rjmp L53: 33000002",
X"addi r1 r14 1: 8b1e0001",
X"cmpi r1 1: e3020001",
X"brne L54: 1f000007",
X"load r0 r14 2 [2]: 810e0002",
X"load r1 r14 24 [2]: 811e0018",
X"mul r0 r0 r1: a7001000",
X"move r2 r0: cf200000",
X"store r14 r2 20 [2]: d1e20014",
X"rjmp L55: 33000005",
X"addi r0 r14 0: 8b0e0000",
X"addi r1 r14 0: 8b1e0000",
X"store r14 r0 20 [2]: d1e00014",
X"store r14 r1 24 [2]: d1e10018",
X"addi r0 r14 0: 8b0e0000",
X"move r12 r14: cfce0000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 478: 8fdd01de",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"load r0 r14 24 [2]: 810e0018",
X"subi r0 r0 1: 8f000001",
X"move r1 r0: cf100000",
X"store r14 r1 24 [2]: d1e10018",
X"cmpi r1 0: e3020000",
X"brge L56: 2f000003",
X"addi r1 r14 0: 8b1e0000",
X"rjmp L57: 33000002",
X"addi r1 r14 1: 8b1e0001",
X"cmpi r1 1: e3020001",
X"brne L58: 1f000007",
X"load r0 r14 2 [2]: 810e0002",
X"load r1 r14 24 [2]: 811e0018",
X"mul r0 r0 r1: a7001000",
X"move r2 r0: cf200000",
X"store r14 r2 20 [2]: d1e20014",
X"rjmp L59: 33000008",
X"load r0 r14 6 [2]: 810e0006",
X"subi r0 r0 1: 8f000001",
X"move r1 r0: cf100000",
X"load r2 r14 4 [2]: 812e0004",
X"move r3 r2: cf320000",
X"store r14 r1 20 [2]: d1e10014",
X"store r14 r3 24 [2]: d1e30018",
X"addi r0 r14 0: 8b0e0000",
X"move r12 r14: cfce0000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 509: 8fdd01fd",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"load r0 r13 2 [1]: 800d0002",
X"load r1 r13 3 [1]: 801d0003",
X"load r2 r14 18 [1]: 802e0012",
X"load r3 r14 10 [2]: 813e000a",
X"cmp r2 r3: df046000",
X"brge L60: 2f000003",
X"addi r2 r14 0: 8b2e0000",
X"rjmp L61: 33000002",
X"addi r2 r14 1: 8b2e0001",
X"load r4 r14 19 [1]: 804e0013",
X"cmp r4 r3: df086000",
X"brge L62: 2f000003",
X"addi r4 r14 0: 8b4e0000",
X"rjmp L63: 33000002",
X"addi r4 r14 1: 8b4e0001",
X"or r2 r2 r4: c3224000",
X"cmpi r2 1: e3040001",
X"brne L64: 1f000007",
X"addi r12 r14 0: 8bce0000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 533: 8fdd0215",
X"rjmprg r13: efd00000",
X"rjmp L65: 33000001",
X"subi r15 r15 2: 8fff0002",
X"load r0 r14 18 [1]: 800e0012",
X"store r13 r0 -2 [2]: d1d0fffe",
X"load r1 r14 19 [1]: 801e0013",
X"add r0 r0 r1: 93001000",
X"move r2 r0: cf200000",
X"subi r15 r15 2: 8fff0002",
X"load r3 r13 2 [1]: 803d0002",
X"store r13 r3 -4 [2]: d1d3fffc",
X"add r3 r3 r2: 93332000",
X"move r4 r3: cf430000",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r5 r13 3 [1]: 805d0003",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r5 0 [2]: d1f50000",
X"subi r15 r15 2: 8fff0002",
X"addi r15 r15 -4: 8bfffffc",
X"store r15 r4 0 [4]: d3f40000",
X"store r13 r2 -2 [2]: d1d2fffe",
X"store r13 r4 -4 [2]: d1d4fffc",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 562: f7d00232",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp tile_index_write: 3300fe2f",
X"addi r15 r15 12: 8bff000c",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r15 r15 4: 8bff0004",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 569: 8fdd0239",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"load r0 r13 2 [1]: 800d0002",
X"load r1 r13 3 [1]: 801d0003",
X"load r2 r13 4 [1]: 802d0004",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r3 r14 2 [2]: 813e0002",
X"add r1 r1 r3: 93113000",
X"mul r1 r1 r2: a7112000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r1 0 [1]: d0f10000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"movlo r13 588: f7d0024c",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp print_c_at: 3300ffb3",
X"addi r15 r15 4: 8bff0004",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 594: 8fdd0252",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"load r0 r13 2 [1]: 800d0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r1 r14 20 [2]: 811e0014",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r1 0 [1]: d0f10000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"movlo r13 609: f7d00261",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp print_c_at: 3300ff9e",
X"addi r15 r15 4: 8bff0004",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"cmpi r12 1: e3180001",
X"brne L66: 1f000016",
X"load r0 r14 20 [2]: 810e0014",
X"addi r0 r0 1: 8b000001",
X"move r1 r0: cf100000",
X"store r14 r1 20 [2]: d1e10014",
X"load r2 r14 6 [2]: 812e0006",
X"cmp r1 r2: df024000",
X"brge L68: 2f000003",
X"addi r1 r14 0: 8b1e0000",
X"rjmp L69: 33000002",
X"addi r1 r14 1: 8b1e0001",
X"cmpi r1 1: e3020001",
X"brne L70: 1f000004",
X"addi r0 r14 0: 8b0e0000",
X"store r14 r0 20 [2]: d1e00014",
X"rjmp L71: 33000001",
X"addi r12 r14 1: 8bce0001",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 633: 8fdd0279",
X"rjmprg r13: efd00000",
X"rjmp L67: 33000001",
X"addi r12 r14 0: 8bce0000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 639: 8fdd027f",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"load r0 r13 4 [2]: 810d0004",
X"load r1 r13 6 [2]: 811d0006",
X"subi r15 r15 2: 8fff0002",
X"addi r2 r14 0: 8b2e0000",
X"store r13 r2 -2 [2]: d1d2fffe",
X"load r0 r13 -2 [2]: 810dfffe",
X"load r1 r13 4 [2]: 811d0004",
X"cmp r0 r1: df002000",
X"brlt L74: 23000003",
X"addi r0 r14 0: 8b0e0000",
X"rjmp L75: 33000002",
X"addi r0 r14 1: 8b0e0001",
X"cmpi r0 1: e3000001",
X"brne L73: 1f000008",
X"load r2 r13 6 [2]: 812d0006",
X"addi r2 r2 1: 8b220001",
X"move r3 r2: cf320000",
X"load r4 r13 -2 [2]: 814dfffe",
X"addi r4 r4 1: 8b440001",
X"move r5 r4: cf540000",
X"rjmp L72: 3300fff1",
X"addi r15 r15 2: 8bff0002",
X"move r12 r14: cfce0000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 667: 8fdd029b",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"subi r15 r15 2: 8fff0002",
X"addi r0 r14 0: 8b0e0000",
X"store r13 r0 -2 [2]: d1d0fffe",
X"load r0 r13 -2 [2]: 810dfffe",
X"load r1 r14 6 [2]: 811e0006",
X"cmp r0 r1: df002000",
X"brlt L78: 23000003",
X"addi r0 r14 0: 8b0e0000",
X"rjmp L79: 33000002",
X"addi r0 r14 1: 8b0e0001",
X"cmpi r0 1: e3000001",
X"brne L77: 1f000013",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"load r2 r13 -2 [2]: 812dfffe",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r2 0 [2]: d1f20000",
X"addi r3 r14 0: 8b3e0000",
X"subi r15 r15 2: 8fff0002",
X"addi r15 r15 -4: 8bfffffc",
X"store r15 r3 0 [4]: d3f30000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 695: f7d002b7",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp tile_index_write: 3300fdaa",
X"addi r15 r15 10: 8bff000a",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"rjmp L76: 3300ffe6",
X"addi r0 r14 0: 8b0e0000",
X"addi r15 r15 2: 8bff0002",
X"move r12 r14: cfce0000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 705: 8fdd02c1",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r0 r14 26 [1]: 800e001a",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r1 r14 0: 8b1e0000",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r1 0 [2]: d1f10000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 723: f7d002d3",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp palette_index_write: 3300fdec",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r0 r14 27 [1]: 800e001b",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r1 r14 1: 8b1e0001",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r1 0 [2]: d1f10000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 742: f7d002e6",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp palette_index_write: 3300fdd9",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r0 r14 28 [1]: 800e001c",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r1 r14 2: 8b1e0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r1 0 [2]: d1f10000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 761: f7d002f9",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp palette_index_write: 3300fdc6",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r0 r14 29 [1]: 800e001d",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r1 r14 3: 8b1e0003",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r1 0 [2]: d1f10000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 780: f7d0030c",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp palette_index_write: 3300fdb3",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r0 r14 30 [1]: 800e001e",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r1 r14 4: 8b1e0004",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r1 0 [2]: d1f10000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 799: f7d0031f",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp palette_index_write: 3300fda0",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r0 r14 31 [1]: 800e001f",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r1 r14 5: 8b1e0005",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r1 0 [2]: d1f10000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 818: f7d00332",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp palette_index_write: 3300fd8d",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r0 r14 32 [1]: 800e0020",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r1 r14 6: 8b1e0006",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r1 0 [2]: d1f10000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 837: f7d00345",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp palette_index_write: 3300fd7a",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r0 r14 33 [1]: 800e0021",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r1 r14 7: 8b1e0007",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r1 0 [2]: d1f10000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 856: f7d00358",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp palette_index_write: 3300fd67",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r0 r14 34 [1]: 800e0022",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r1 r14 8: 8b1e0008",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r1 0 [2]: d1f10000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 875: f7d0036b",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp palette_index_write: 3300fd54",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r0 r14 35 [1]: 800e0023",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r1 r14 9: 8b1e0009",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r1 0 [2]: d1f10000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 894: f7d0037e",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp palette_index_write: 3300fd41",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r0 r14 36 [1]: 800e0024",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r1 r14 10: 8b1e000a",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r1 0 [2]: d1f10000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 913: f7d00391",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp palette_index_write: 3300fd2e",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r0 r14 37 [1]: 800e0025",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r1 r14 11: 8b1e000b",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r1 0 [2]: d1f10000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 932: f7d003a4",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp palette_index_write: 3300fd1b",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r0 r14 38 [1]: 800e0026",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r1 r14 12: 8b1e000c",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r1 0 [2]: d1f10000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 951: f7d003b7",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp palette_index_write: 3300fd08",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r0 r14 39 [1]: 800e0027",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r1 r14 13: 8b1e000d",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r1 0 [2]: d1f10000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 970: f7d003ca",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp palette_index_write: 3300fcf5",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"load r0 r14 40 [1]: 800e0028",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r1 r14 14: 8b1e000e",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r1 0 [2]: d1f10000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 989: f7d003dd",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp palette_index_write: 3300fce2",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"addi r0 r14 0: 8b0e0000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r0 r14 0: 8b0e0000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r0 0 [1]: d0f00000",
X"addi r0 r14 15: 8b0e000f",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r0 0 [2]: d1f00000",
X"subi r15 r15 2: 8fff0002",
X"movlo r13 1009: f7d003f1",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp palette_index_write: 3300fcce",
X"addi r15 r15 8: 8bff0008",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"move r12 r14: cfce0000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 1016: 8fdd03f8",
X"rjmprg r13: efd00000",
X"move r13 r15: cfdf0000",
X"subi r15 r15 2: 8fff0002",
X"addi r0 r14 0: 8b0e0000",
X"subi r15 r15 2: 8fff0002",
X"addi r1 r14 0: 8b1e0000",
X"store r13 r0 -2 [2]: d1d0fffe",
X"store r13 r1 -4 [2]: d1d1fffc",
X"load r0 r13 -2 [2]: 810dfffe",
X"load r1 r14 6 [2]: 811e0006",
X"cmp r0 r1: df002000",
X"brlt L82: 23000003",
X"addi r0 r14 0: 8b0e0000",
X"rjmp L83: 33000002",
X"addi r0 r14 1: 8b0e0001",
X"cmpi r0 1: e3000001",
X"brne L81: 1f000025",
X"load r2 r13 -4 [2]: 812dfffc",
X"cmpi r2 11: e304000b",
X"brge L84: 2f000003",
X"addi r2 r14 0: 8b2e0000",
X"rjmp L85: 33000002",
X"addi r2 r14 1: 8b2e0001",
X"cmpi r2 1: e3040001",
X"brne L86: 1f000004",
X"addi r0 r14 0: 8b0e0000",
X"store r13 r0 -4 [2]: d1d0fffc",
X"rjmp L87: 33000001",
X"addi r0 r14 4: 8b0e0004",
X"load r1 r13 -4 [2]: 811dfffc",
X"add r0 r0 r1: 93001000",
X"move r2 r0: cf200000",
X"addi r15 r15 -2: 8bfffffe",
X"store r15 r13 0 [2]: d1fd0000",
X"subi r15 r15 2: 8fff0002",
X"addi r3 r14 0: 8b3e0000",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r3 0 [1]: d0f30000",
X"store r14 r2 19 [1]: d0e20013",
X"movlo r13 1059: f7d00423",
X"addi r15 r15 -1: 8bffffff",
X"store r15 r13 0: d3fd0000",
X"rjmp print_c: 3300fe31",
X"addi r15 r15 3: 8bff0003",
X"load r13 r15 0 [2]: 81df0000",
X"addi r15 r15 2: 8bff0002",
X"load r0 r13 -2 [2]: 810dfffe",
X"addi r0 r0 1: 8b000001",
X"move r1 r0: cf100000",
X"load r2 r13 -4 [2]: 812dfffc",
X"addi r2 r2 1: 8b220001",
X"move r3 r2: cf320000",
X"rjmp L80: 3300ffd4",
X"addi r15 r15 4: 8bff0004",
X"move r12 r14: cfce0000",
X"load r13 r15 0: 83df0000",
X"addi r15 r15 1: 8bff0001",
X"subi r13 r13 1074: 8fdd0432",
X"rjmprg r13: efd00000",
--$PROGRAM_END
others => X"00000000"
);