mem := (
--$DATA

--$DATA_END
)