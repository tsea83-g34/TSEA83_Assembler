mem := (
--$PROGRAM
"00110011000000000000000000001111",
"10001111011001100000000000000001",
"11010011011000000000001000000000",
"00110011000000000000000000001100",
"111000110001011000000000001000000",
"00011011000000001111111111111100",
"110100110110101100000010000000000",
"1000111110101010000000000000100000",
"10001011011001100000000000000001",
"00110011000000000000000000000110",
"00111111000100000000000000001000",
"101111110001101000010000000000000",
"11100011000000100000000000000001",
"00100111000000001111111111110111",
"00110011000000000000000000000001",
"00110011000000001111111111111011",
--$PROGRAM_END
others => X"00000000"
);