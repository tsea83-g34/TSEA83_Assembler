mem := (
--$PROGRAM
X"93001000",
X"8b110001",
X"83df0000",
X"8bff0001",
X"8fdd0005",
X"efd00000",
X"f7d0000a",
X"d3fd0000",
X"8bffffff",
X"3300fff8",
--$PROGRAM_END
others => X"00000000"
);