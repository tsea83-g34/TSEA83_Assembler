mem := (
--$PROGRAM
X"07000011",
X"07100000",
X"07200000",
X"471e0004",
X"472e0003",
X"cf024000",
X"0b000006",
X"131f0000",
X"07200000",
X"07100000",
X"07f00000",
X"1f000000",
X"132f0000",
X"07200000",
X"07100000",
X"07f00000",
X"1f000000",
X"171a000a",
X"2e540028",
X"07100000",
X"07200000",
X"1f00ffec",
X"07300000"
--$PROGRAM_END
);