library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library work;
use work.PIPECPU_STD.ALL;

package program_file is
  
  constant program : program_memory_array := (
--$PROGRAM
"10001011000100010000000000000001", -- addi r1 r1 1
"10001011001000100000000000000010", -- addi r2 r2 2
"10001011001100110000000000000011", -- addi r3 r3 3
"11010011001100110000000000000000", -- store r3 r3 0 [4]
"10000011010100110000000000000000", -- load r5 r3 0 [4]
"10001011010101010000000000000001", -- addi r5 r5 1 [ADD_r5]
"11100011000001010000000000000101", -- cmpi r5 5
"00011111000000001111111111111110", -- brne ADD_r5
"10001011101010101111111011011100", -- addi r10 r10 0xfedc
"11010001000010100000000000001010", -- store r0 r10 10 [1]
"10000001101000000000000000001010", -- load r10 r0 10 [1]
"11110111110111010000000000001111", -- movlo r13 r13 15
"10001011111111111111111111111110", -- addi r15 r15 -2
"11010010111111010000000000000000", -- store r15 r13 0 [2]
"00110011000000000000000000001101", -- rjmp SUBROUTINE
"00000011000000000000000000000000", -- nop
"00000011000000000000000000000000", -- nop
"00000011000000000000000000000000", -- nop
"00000011000000000000000000000000", -- nop
"00000011000000000000000000000000", -- nop
"00000011000000000000000000000000", -- nop
"00000011000000000000000000000000", -- nop
"00000011000000000000000000000000", -- nop
"00000011000000000000000000000000", -- nop
"00000011000000000000000000000000", -- nop
"00000011000000000000000000000000", -- nop
"00000011000000000000000000000000", -- nop
"10000010110111110000000000000000", -- load r13 r15 0 [2] [SUBROUTINE]
"10001011111111110000000000000010", -- addi r15 r15 2
"10001111110111010000000000011110", -- subi r13 r13 30
"11101111000011010000000000000000", -- rjmprg r13
--$PROGRAM_END
others => X"00000000"
);

end program_file;
