mem := (
--$DATA
X"00",
X"10",
X"28",
X"00",
X"1e",
X"00",
X"00",
X"00",
X"00",
X"00",
X"10",
X"00",
X"00",
X"00",
X"80",
X"02",
X"e0",
X"01",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"00",
X"49",
X"92",
X"ff",
X"e0",
X"f0",
X"fc",
X"9c",
X"1c",
X"1e",
X"1f",
X"13",
X"03",
X"83",
X"e3",
X"5f",
X"fd",
X"be",
X"2d",
X"6c",
X"4d",
X"cf",
X"24",
X"76",
X"b6",
X"57",
X"e9",
--$DATA_END
others => X"00"
)